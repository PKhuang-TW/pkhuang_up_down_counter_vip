`ifndef COUNTER_PACKAGE_SV
`define COUNTER_PACKAGE_SV

package counter_package;
    parameter P_ADDR_WIDTH = 3;
endpackage

`endif